LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY LATCH_ADDR IS
PORT
(
	AD : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
	A16 : IN STD_LOGIC;
	A17 : IN STD_LOGIC;
	A18 : IN STD_LOGIC;
	NADV : IN STD_LOGIC;
	NOE : IN STD_LOGIC;
	NWE : IN STD_LOGIC;
   ADDR : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
	CS0 : OUT STD_LOGIC;
	CS1 : OUT STD_LOGIC;
	CS2 : OUT STD_LOGIC; 
	CS3 : OUT STD_LOGIC;
	CS4 : OUT STD_LOGIC;
	CS5 : OUT STD_LOGIC;
	CS6 : OUT STD_LOGIC;
	CS7 : OUT STD_LOGIC;
	nCS : OUT STD_LOGIC
);
END LATCH_ADDR;

ARCHITECTURE LATCH OF LATCH_ADDR IS
BEGIN
	PROCESS(NADV,AD,A16,A17,A18,NOE,NWE)
	BEGIN
		IF(NADV'EVENT and NADV='1' AND (NWE = '1' OR NOE = '1'))THEN
			ADDR<=AD;
			nCS <= NOT A16;
			IF(A16 = '1') THEN
				IF(AD(15 DOWNTO 8) = X"80") THEN
					CS0<='0';CS1<='1';CS2<='1';CS3<='1';
					CS4<='1';CS5<='1';CS6<='1';CS7<='1';
				ELSIF(AD(15 DOWNTO 8) = X"81") THEN
					CS0<='1';CS1<='0';CS2<='1';CS3<='1';
					CS4<='1';CS5<='1';CS6<='1';CS7<='1';
				ELSIF(AD(15 DOWNTO 8) = X"82") THEN
					CS0<='1';CS1<='1';CS2<='0';CS3<='1';
					CS4<='1';CS5<='1';CS6<='1';CS7<='1';
				ELSIF(AD(15 DOWNTO 8) = X"83") THEN
					CS0<='1';CS1<='1';CS2<='1';CS3<='0';
					CS4<='1';CS5<='1';CS6<='1';CS7<='1';
				ELSIF(AD(15 DOWNTO 8) = X"84") THEN
					CS0<='1';CS1<='1';CS2<='1';CS3<='1';
					CS4<='0';CS5<='1';CS6<='1';CS7<='1';
				ELSIF(AD(15 DOWNTO 8) = X"85") THEN
					CS0<='1';CS1<='1';CS2<='1';CS3<='1';
					CS4<='1';CS5<='0';CS6<='1';CS7<='1';
				ELSIF(AD(15 DOWNTO 8) = X"86") THEN
					CS0<='1';CS1<='1';CS2<='1';CS3<='1';
					CS4<='1';CS5<='1';CS6<='0';CS7<='1';
				ELSIF(AD(15 DOWNTO 8) = X"87") THEN
					CS0<='1';CS1<='1';CS2<='1';CS3<='1';
					CS4<='1';CS5<='1';CS6<='1';CS7<='0';
				ELSE
					CS0<='1';CS1<='1';CS2<='1';CS3<='1';
					CS4<='1';CS5<='1';CS6<='1';CS7<='1';
				END IF;
			ELSE
					CS0<='1';CS1<='1';CS2<='1';CS3<='1';
					CS4<='1';CS5<='1';CS6<='1';CS7<='1';
			END IF;
		END IF;
	END PROCESS;
END LATCH;