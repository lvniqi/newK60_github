LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY DECODER_ADDR IS
PORT
(
	ADDR : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
	CS0 : IN STD_LOGIC;
	CS_FREQ_WR_L : OUT STD_LOGIC;
	CS_FREQ_WR_H : OUT STD_LOGIC;
	CS_FREQ_RD_L : OUT STD_LOGIC;
	CS_FREQ_RD_H : OUT STD_LOGIC
);
END DECODER_ADDR;

ARCHITECTURE DECODER OF DECODER_ADDR IS
BEGIN
	PROCESS(CS0, ADDR)
	BEGIN
		IF(CS0 = '0')THEN
			IF(ADDR(7 DOWNTO 0)=X"00")THEN
				CS_FREQ_WR_L<='0';CS_FREQ_WR_H<='1';
				CS_FREQ_RD_L<='1';CS_FREQ_RD_H<='1';
			ELSIF(ADDR(7 DOWNTO 0)=X"01")THEN
				CS_FREQ_WR_L<='1';CS_FREQ_WR_H<='0';
				CS_FREQ_RD_L<='1';CS_FREQ_RD_H<='1';
			ELSIF(ADDR(7 DOWNTO 0)=X"02")THEN
				CS_FREQ_WR_L<='1';CS_FREQ_WR_H<='1';
				CS_FREQ_RD_L<='0';CS_FREQ_RD_H<='1';
			ELSIF(ADDR(7 DOWNTO 0)=X"03")THEN
				CS_FREQ_WR_L<='1';CS_FREQ_WR_H<='1';
				CS_FREQ_RD_L<='1';CS_FREQ_RD_H<='0';
			ELSE
				CS_FREQ_WR_L<='1';CS_FREQ_WR_H<='1';
				CS_FREQ_RD_L<='1';CS_FREQ_RD_H<='1';
			END IF;
		ELSE
			CS_FREQ_WR_L<='1';CS_FREQ_WR_H<='1';
			CS_FREQ_RD_L<='1';CS_FREQ_RD_H<='1';
		END IF;
	END PROCESS;	
END DECODER;