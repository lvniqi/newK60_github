LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY LATCH_AD IS
PORT
(
	AD : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
   DATA : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
   NADV : IN STD_LOGIC;
	NOE : IN STD_LOGIC;
	NWE : IN STD_LOGIC;
	nCS : IN STD_LOGIC
);
END LATCH_AD;

ARCHITECTURE D2AD OF LATCH_AD IS
BEGIN
	PROCESS(NWE,NOE,nCS,DATA)
	BEGIN
		IF(nCS='0')THEN
			IF( NWE = '1' AND NOE='0' AND NADV = '1')THEN
				AD<=DATA;
			ELSE
				AD<=(OTHERS=>'Z');
			END IF;
		ELSE 
			AD<=(OTHERS=>'Z');
		END IF;
	END PROCESS;
END D2AD;