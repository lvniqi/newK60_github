LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY LATCH_DATA IS
    PORT(
	 NADV : In STD_LOGIC;
        AD : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
        DATA : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
        NOE : In STD_LOGIC;
		NWE : IN STD_LOGIC;
		nCS : IN STD_LOGIC
		);
END LATCH_DATA;

ARCHITECTURE AD2D OF LATCH_DATA IS
BEGIN
	PROCESS(NWE,NOE,nCS,AD)
	BEGIN
		IF(nCS='0')THEN
			IF( NWE='0'AND NOE='1' AND NADV = '1')THEN
			--DATA<="0000000000000110";
				DATA<=AD;
			ELSIF(NOE='0')THEN
				DATA<=(OTHERS=>'Z');
			END IF;
		ELSE 
			DATA<=(OTHERS=>'Z');
		END IF;
	END PROCESS;
END AD2D;